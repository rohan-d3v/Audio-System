/*
Rohan Krishna Ramkhumar, rxr353
Sydney Tenaglia, snt21
*/
module digital(
					input clk,
					input din,
					output dout,
					output [11:0] res,
					output cs,
					output valid
					);