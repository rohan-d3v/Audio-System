/*
Rohan Krishna Ramkhumar, rxr353
Sydney Tenaglia, snt21
*/

module peakrst()